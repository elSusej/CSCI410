module bit_test;
  reg in, load;
  wire out;

  student_bit dut (.in(in), .load(load), .out(out));

  initial begin
    $display("|time|in|load|out|");

    in = 1'b0;
    load = 1'b0;
    #1 $display("|0+|%b|%b|%b|", in, load, out);

    in = 1'b0;
    load = 1'b0;
    #1 $display("|1|%b|%b|%b|", in, load, out);

    in = 1'b0;
    load = 1'b1;
    #1 $display("|1+|%b|%b|%b|", in, load, out);

    in = 1'b0;
    load = 1'b1;
    #1 $display("|2|%b|%b|%b|", in, load, out);

    in = 1'b1;
    load = 1'b0;
    #1 $display("|2+|%b|%b|%b|", in, load, out);

    in = 1'b1;
    load = 1'b0;
    #1 $display("|3|%b|%b|%b|", in, load, out);

    in = 1'b1;
    load = 1'b1;
    #1 $display("|3+|%b|%b|%b|", in, load, out);

    in = 1'b1;
    load = 1'b1;
    #1 $display("|4|%b|%b|%b|", in, load, out);

    in = 1'b0;
    load = 1'b0;
    #1 $display("|4+|%b|%b|%b|", in, load, out);

    in = 1'b0;
    load = 1'b0;
    #1 $display("|5|%b|%b|%b|", in, load, out);

    in = 1'b1;
    load = 1'b0;
    #1 $display("|5+|%b|%b|%b|", in, load, out);

    in = 1'b1;
    load = 1'b0;
    #1 $display("|6|%b|%b|%b|", in, load, out);

    in = 1'b0;
    load = 1'b1;
    #1 $display("|6+|%b|%b|%b|", in, load, out);

    in = 1'b0;
    load = 1'b1;
    #1 $display("|7|%b|%b|%b|", in, load, out);

    in = 1'b1;
    load = 1'b1;
    #1 $display("|7+|%b|%b|%b|", in, load, out);

    in = 1'b1;
    load = 1'b1;
    #1 $display("|8|%b|%b|%b|", in, load, out);

    in = 1'b0;
    load = 1'b0;
    #1 $display("|8+|%b|%b|%b|", in, load, out);

    in = 1'b0;
    load = 1'b0;
    #1 $display("|9|%b|%b|%b|", in, load, out);

    in = 1'b0;
    load = 1'b0;
    #1 $display("|9+|%b|%b|%b|", in, load, out);

    in = 1'b0;
    load = 1'b0;
    #1 $display("|10|%b|%b|%b|", in, load, out);

    in = 1'b0;
    load = 1'b0;
    #1 $display("|10+|%b|%b|%b|", in, load, out);

    in = 1'b0;
    load = 1'b0;
    #1 $display("|11|%b|%b|%b|", in, load, out);

    in = 1'b0;
    load = 1'b0;
    #1 $display("|11+|%b|%b|%b|", in, load, out);

    in = 1'b0;
    load = 1'b0;
    #1 $display("|12|%b|%b|%b|", in, load, out);

    in = 1'b0;
    load = 1'b0;
    #1 $display("|12+|%b|%b|%b|", in, load, out);

    in = 1'b0;
    load = 1'b0;
    #1 $display("|13|%b|%b|%b|", in, load, out);

    in = 1'b0;
    load = 1'b0;
    #1 $display("|13+|%b|%b|%b|", in, load, out);

    in = 1'b0;
    load = 1'b0;
    #1 $display("|14|%b|%b|%b|", in, load, out);

    in = 1'b0;
    load = 1'b0;
    #1 $display("|14+|%b|%b|%b|", in, load, out);

    in = 1'b0;
    load = 1'b0;
    #1 $display("|15|%b|%b|%b|", in, load, out);

    in = 1'b0;
    load = 1'b0;
    #1 $display("|15+|%b|%b|%b|", in, load, out);

    in = 1'b0;
    load = 1'b0;
    #1 $display("|16|%b|%b|%b|", in, load, out);

    in = 1'b0;
    load = 1'b0;
    #1 $display("|16+|%b|%b|%b|", in, load, out);

    in = 1'b0;
    load = 1'b0;
    #1 $display("|17|%b|%b|%b|", in, load, out);

    in = 1'b0;
    load = 1'b0;
    #1 $display("|17+|%b|%b|%b|", in, load, out);

    in = 1'b0;
    load = 1'b0;
    #1 $display("|18|%b|%b|%b|", in, load, out);

    in = 1'b0;
    load = 1'b0;
    #1 $display("|18+|%b|%b|%b|", in, load, out);

    in = 1'b0;
    load = 1'b0;
    #1 $display("|19|%b|%b|%b|", in, load, out);

    in = 1'b0;
    load = 1'b0;
    #1 $display("|19+|%b|%b|%b|", in, load, out);

    in = 1'b0;
    load = 1'b0;
    #1 $display("|20|%b|%b|%b|", in, load, out);

    in = 1'b0;
    load = 1'b0;
    #1 $display("|20+|%b|%b|%b|", in, load, out);

    in = 1'b0;
    load = 1'b0;
    #1 $display("|21|%b|%b|%b|", in, load, out);

    in = 1'b0;
    load = 1'b0;
    #1 $display("|21+|%b|%b|%b|", in, load, out);

    in = 1'b0;
    load = 1'b0;
    #1 $display("|22|%b|%b|%b|", in, load, out);

    in = 1'b0;
    load = 1'b0;
    #1 $display("|22+|%b|%b|%b|", in, load, out);

    in = 1'b0;
    load = 1'b0;
    #1 $display("|23|%b|%b|%b|", in, load, out);

    in = 1'b0;
    load = 1'b0;
    #1 $display("|23+|%b|%b|%b|", in, load, out);

    in = 1'b0;
    load = 1'b0;
    #1 $display("|24|%b|%b|%b|", in, load, out);

    in = 1'b0;
    load = 1'b0;
    #1 $display("|24+|%b|%b|%b|", in, load, out);

    in = 1'b0;
    load = 1'b0;
    #1 $display("|25|%b|%b|%b|", in, load, out);

    in = 1'b0;
    load = 1'b0;
    #1 $display("|25+|%b|%b|%b|", in, load, out);

    in = 1'b0;
    load = 1'b0;
    #1 $display("|26|%b|%b|%b|", in, load, out);

    in = 1'b0;
    load = 1'b0;
    #1 $display("|26+|%b|%b|%b|", in, load, out);

    in = 1'b0;
    load = 1'b0;
    #1 $display("|27|%b|%b|%b|", in, load, out);

    in = 1'b0;
    load = 1'b0;
    #1 $display("|27+|%b|%b|%b|", in, load, out);

    in = 1'b0;
    load = 1'b0;
    #1 $display("|28|%b|%b|%b|", in, load, out);

    in = 1'b0;
    load = 1'b0;
    #1 $display("|28+|%b|%b|%b|", in, load, out);

    in = 1'b0;
    load = 1'b0;
    #1 $display("|29|%b|%b|%b|", in, load, out);

    in = 1'b0;
    load = 1'b0;
    #1 $display("|29+|%b|%b|%b|", in, load, out);

    in = 1'b0;
    load = 1'b0;
    #1 $display("|30|%b|%b|%b|", in, load, out);

    in = 1'b0;
    load = 1'b0;
    #1 $display("|30+|%b|%b|%b|", in, load, out);

    in = 1'b0;
    load = 1'b0;
    #1 $display("|31|%b|%b|%b|", in, load, out);

    in = 1'b0;
    load = 1'b0;
    #1 $display("|31+|%b|%b|%b|", in, load, out);

    in = 1'b0;
    load = 1'b0;
    #1 $display("|32|%b|%b|%b|", in, load, out);

    in = 1'b0;
    load = 1'b0;
    #1 $display("|32+|%b|%b|%b|", in, load, out);

    in = 1'b0;
    load = 1'b0;
    #1 $display("|33|%b|%b|%b|", in, load, out);

    in = 1'b0;
    load = 1'b0;
    #1 $display("|33+|%b|%b|%b|", in, load, out);

    in = 1'b0;
    load = 1'b0;
    #1 $display("|34|%b|%b|%b|", in, load, out);

    in = 1'b0;
    load = 1'b0;
    #1 $display("|34+|%b|%b|%b|", in, load, out);

    in = 1'b0;
    load = 1'b0;
    #1 $display("|35|%b|%b|%b|", in, load, out);

    in = 1'b0;
    load = 1'b0;
    #1 $display("|35+|%b|%b|%b|", in, load, out);

    in = 1'b0;
    load = 1'b0;
    #1 $display("|36|%b|%b|%b|", in, load, out);

    in = 1'b0;
    load = 1'b0;
    #1 $display("|36+|%b|%b|%b|", in, load, out);

    in = 1'b0;
    load = 1'b0;
    #1 $display("|37|%b|%b|%b|", in, load, out);

    in = 1'b0;
    load = 1'b0;
    #1 $display("|37+|%b|%b|%b|", in, load, out);

    in = 1'b0;
    load = 1'b0;
    #1 $display("|38|%b|%b|%b|", in, load, out);

    in = 1'b0;
    load = 1'b0;
    #1 $display("|38+|%b|%b|%b|", in, load, out);

    in = 1'b0;
    load = 1'b0;
    #1 $display("|39|%b|%b|%b|", in, load, out);

    in = 1'b0;
    load = 1'b0;
    #1 $display("|39+|%b|%b|%b|", in, load, out);

    in = 1'b0;
    load = 1'b0;
    #1 $display("|40|%b|%b|%b|", in, load, out);

    in = 1'b0;
    load = 1'b0;
    #1 $display("|40+|%b|%b|%b|", in, load, out);

    in = 1'b0;
    load = 1'b0;
    #1 $display("|41|%b|%b|%b|", in, load, out);

    in = 1'b0;
    load = 1'b0;
    #1 $display("|41+|%b|%b|%b|", in, load, out);

    in = 1'b0;
    load = 1'b0;
    #1 $display("|42|%b|%b|%b|", in, load, out);

    in = 1'b0;
    load = 1'b0;
    #1 $display("|42+|%b|%b|%b|", in, load, out);

    in = 1'b0;
    load = 1'b0;
    #1 $display("|43|%b|%b|%b|", in, load, out);

    in = 1'b0;
    load = 1'b0;
    #1 $display("|43+|%b|%b|%b|", in, load, out);

    in = 1'b0;
    load = 1'b0;
    #1 $display("|44|%b|%b|%b|", in, load, out);

    in = 1'b0;
    load = 1'b0;
    #1 $display("|44+|%b|%b|%b|", in, load, out);

    in = 1'b0;
    load = 1'b0;
    #1 $display("|45|%b|%b|%b|", in, load, out);

    in = 1'b0;
    load = 1'b0;
    #1 $display("|45+|%b|%b|%b|", in, load, out);

    in = 1'b0;
    load = 1'b0;
    #1 $display("|46|%b|%b|%b|", in, load, out);

    in = 1'b0;
    load = 1'b0;
    #1 $display("|46+|%b|%b|%b|", in, load, out);

    in = 1'b0;
    load = 1'b0;
    #1 $display("|47|%b|%b|%b|", in, load, out);

    in = 1'b0;
    load = 1'b0;
    #1 $display("|47+|%b|%b|%b|", in, load, out);

    in = 1'b0;
    load = 1'b0;
    #1 $display("|48|%b|%b|%b|", in, load, out);

    in = 1'b0;
    load = 1'b0;
    #1 $display("|48+|%b|%b|%b|", in, load, out);

    in = 1'b0;
    load = 1'b0;
    #1 $display("|49|%b|%b|%b|", in, load, out);

    in = 1'b0;
    load = 1'b0;
    #1 $display("|49+|%b|%b|%b|", in, load, out);

    in = 1'b0;
    load = 1'b0;
    #1 $display("|50|%b|%b|%b|", in, load, out);

    in = 1'b0;
    load = 1'b0;
    #1 $display("|50+|%b|%b|%b|", in, load, out);

    in = 1'b0;
    load = 1'b0;
    #1 $display("|51|%b|%b|%b|", in, load, out);

    in = 1'b0;
    load = 1'b0;
    #1 $display("|51+|%b|%b|%b|", in, load, out);

    in = 1'b0;
    load = 1'b0;
    #1 $display("|52|%b|%b|%b|", in, load, out);

    in = 1'b0;
    load = 1'b0;
    #1 $display("|52+|%b|%b|%b|", in, load, out);

    in = 1'b0;
    load = 1'b0;
    #1 $display("|53|%b|%b|%b|", in, load, out);

    in = 1'b0;
    load = 1'b0;
    #1 $display("|53+|%b|%b|%b|", in, load, out);

    in = 1'b0;
    load = 1'b0;
    #1 $display("|54|%b|%b|%b|", in, load, out);

    in = 1'b0;
    load = 1'b0;
    #1 $display("|54+|%b|%b|%b|", in, load, out);

    in = 1'b0;
    load = 1'b0;
    #1 $display("|55|%b|%b|%b|", in, load, out);

    in = 1'b0;
    load = 1'b0;
    #1 $display("|55+|%b|%b|%b|", in, load, out);

    in = 1'b0;
    load = 1'b0;
    #1 $display("|56|%b|%b|%b|", in, load, out);

    in = 1'b0;
    load = 1'b0;
    #1 $display("|56+|%b|%b|%b|", in, load, out);

    in = 1'b0;
    load = 1'b0;
    #1 $display("|57|%b|%b|%b|", in, load, out);

    in = 1'b0;
    load = 1'b1;
    #1 $display("|57+|%b|%b|%b|", in, load, out);

    in = 1'b0;
    load = 1'b1;
    #1 $display("|58|%b|%b|%b|", in, load, out);

    in = 1'b1;
    load = 1'b0;
    #1 $display("|58+|%b|%b|%b|", in, load, out);

    in = 1'b1;
    load = 1'b0;
    #1 $display("|59|%b|%b|%b|", in, load, out);

    in = 1'b1;
    load = 1'b0;
    #1 $display("|59+|%b|%b|%b|", in, load, out);

    in = 1'b1;
    load = 1'b0;
    #1 $display("|60|%b|%b|%b|", in, load, out);

    in = 1'b1;
    load = 1'b0;
    #1 $display("|60+|%b|%b|%b|", in, load, out);

    in = 1'b1;
    load = 1'b0;
    #1 $display("|61|%b|%b|%b|", in, load, out);

    in = 1'b1;
    load = 1'b0;
    #1 $display("|61+|%b|%b|%b|", in, load, out);

    in = 1'b1;
    load = 1'b0;
    #1 $display("|62|%b|%b|%b|", in, load, out);

    in = 1'b1;
    load = 1'b0;
    #1 $display("|62+|%b|%b|%b|", in, load, out);

    in = 1'b1;
    load = 1'b0;
    #1 $display("|63|%b|%b|%b|", in, load, out);

    in = 1'b1;
    load = 1'b0;
    #1 $display("|63+|%b|%b|%b|", in, load, out);

    in = 1'b1;
    load = 1'b0;
    #1 $display("|64|%b|%b|%b|", in, load, out);

    in = 1'b1;
    load = 1'b0;
    #1 $display("|64+|%b|%b|%b|", in, load, out);

    in = 1'b1;
    load = 1'b0;
    #1 $display("|65|%b|%b|%b|", in, load, out);

    in = 1'b1;
    load = 1'b0;
    #1 $display("|65+|%b|%b|%b|", in, load, out);

    in = 1'b1;
    load = 1'b0;
    #1 $display("|66|%b|%b|%b|", in, load, out);

    in = 1'b1;
    load = 1'b0;
    #1 $display("|66+|%b|%b|%b|", in, load, out);

    in = 1'b1;
    load = 1'b0;
    #1 $display("|67|%b|%b|%b|", in, load, out);

    in = 1'b1;
    load = 1'b0;
    #1 $display("|67+|%b|%b|%b|", in, load, out);

    in = 1'b1;
    load = 1'b0;
    #1 $display("|68|%b|%b|%b|", in, load, out);

    in = 1'b1;
    load = 1'b0;
    #1 $display("|68+|%b|%b|%b|", in, load, out);

    in = 1'b1;
    load = 1'b0;
    #1 $display("|69|%b|%b|%b|", in, load, out);

    in = 1'b1;
    load = 1'b0;
    #1 $display("|69+|%b|%b|%b|", in, load, out);

    in = 1'b1;
    load = 1'b0;
    #1 $display("|70|%b|%b|%b|", in, load, out);

    in = 1'b1;
    load = 1'b0;
    #1 $display("|70+|%b|%b|%b|", in, load, out);

    in = 1'b1;
    load = 1'b0;
    #1 $display("|71|%b|%b|%b|", in, load, out);

    in = 1'b1;
    load = 1'b0;
    #1 $display("|71+|%b|%b|%b|", in, load, out);

    in = 1'b1;
    load = 1'b0;
    #1 $display("|72|%b|%b|%b|", in, load, out);

    in = 1'b1;
    load = 1'b0;
    #1 $display("|72+|%b|%b|%b|", in, load, out);

    in = 1'b1;
    load = 1'b0;
    #1 $display("|73|%b|%b|%b|", in, load, out);

    in = 1'b1;
    load = 1'b0;
    #1 $display("|73+|%b|%b|%b|", in, load, out);

    in = 1'b1;
    load = 1'b0;
    #1 $display("|74|%b|%b|%b|", in, load, out);

    in = 1'b1;
    load = 1'b0;
    #1 $display("|74+|%b|%b|%b|", in, load, out);

    in = 1'b1;
    load = 1'b0;
    #1 $display("|75|%b|%b|%b|", in, load, out);

    in = 1'b1;
    load = 1'b0;
    #1 $display("|75+|%b|%b|%b|", in, load, out);

    in = 1'b1;
    load = 1'b0;
    #1 $display("|76|%b|%b|%b|", in, load, out);

    in = 1'b1;
    load = 1'b0;
    #1 $display("|76+|%b|%b|%b|", in, load, out);

    in = 1'b1;
    load = 1'b0;
    #1 $display("|77|%b|%b|%b|", in, load, out);

    in = 1'b1;
    load = 1'b0;
    #1 $display("|77+|%b|%b|%b|", in, load, out);

    in = 1'b1;
    load = 1'b0;
    #1 $display("|78|%b|%b|%b|", in, load, out);

    in = 1'b1;
    load = 1'b0;
    #1 $display("|78+|%b|%b|%b|", in, load, out);

    in = 1'b1;
    load = 1'b0;
    #1 $display("|79|%b|%b|%b|", in, load, out);

    in = 1'b1;
    load = 1'b0;
    #1 $display("|79+|%b|%b|%b|", in, load, out);

    in = 1'b1;
    load = 1'b0;
    #1 $display("|80|%b|%b|%b|", in, load, out);

    in = 1'b1;
    load = 1'b0;
    #1 $display("|80+|%b|%b|%b|", in, load, out);

    in = 1'b1;
    load = 1'b0;
    #1 $display("|81|%b|%b|%b|", in, load, out);

    in = 1'b1;
    load = 1'b0;
    #1 $display("|81+|%b|%b|%b|", in, load, out);

    in = 1'b1;
    load = 1'b0;
    #1 $display("|82|%b|%b|%b|", in, load, out);

    in = 1'b1;
    load = 1'b0;
    #1 $display("|82+|%b|%b|%b|", in, load, out);

    in = 1'b1;
    load = 1'b0;
    #1 $display("|83|%b|%b|%b|", in, load, out);

    in = 1'b1;
    load = 1'b0;
    #1 $display("|83+|%b|%b|%b|", in, load, out);

    in = 1'b1;
    load = 1'b0;
    #1 $display("|84|%b|%b|%b|", in, load, out);

    in = 1'b1;
    load = 1'b0;
    #1 $display("|84+|%b|%b|%b|", in, load, out);

    in = 1'b1;
    load = 1'b0;
    #1 $display("|85|%b|%b|%b|", in, load, out);

    in = 1'b1;
    load = 1'b0;
    #1 $display("|85+|%b|%b|%b|", in, load, out);

    in = 1'b1;
    load = 1'b0;
    #1 $display("|86|%b|%b|%b|", in, load, out);

    in = 1'b1;
    load = 1'b0;
    #1 $display("|86+|%b|%b|%b|", in, load, out);

    in = 1'b1;
    load = 1'b0;
    #1 $display("|87|%b|%b|%b|", in, load, out);

    in = 1'b1;
    load = 1'b0;
    #1 $display("|87+|%b|%b|%b|", in, load, out);

    in = 1'b1;
    load = 1'b0;
    #1 $display("|88|%b|%b|%b|", in, load, out);

    in = 1'b1;
    load = 1'b0;
    #1 $display("|88+|%b|%b|%b|", in, load, out);

    in = 1'b1;
    load = 1'b0;
    #1 $display("|89|%b|%b|%b|", in, load, out);

    in = 1'b1;
    load = 1'b0;
    #1 $display("|89+|%b|%b|%b|", in, load, out);

    in = 1'b1;
    load = 1'b0;
    #1 $display("|90|%b|%b|%b|", in, load, out);

    in = 1'b1;
    load = 1'b0;
    #1 $display("|90+|%b|%b|%b|", in, load, out);

    in = 1'b1;
    load = 1'b0;
    #1 $display("|91|%b|%b|%b|", in, load, out);

    in = 1'b1;
    load = 1'b0;
    #1 $display("|91+|%b|%b|%b|", in, load, out);

    in = 1'b1;
    load = 1'b0;
    #1 $display("|92|%b|%b|%b|", in, load, out);

    in = 1'b1;
    load = 1'b0;
    #1 $display("|92+|%b|%b|%b|", in, load, out);

    in = 1'b1;
    load = 1'b0;
    #1 $display("|93|%b|%b|%b|", in, load, out);

    in = 1'b1;
    load = 1'b0;
    #1 $display("|93+|%b|%b|%b|", in, load, out);

    in = 1'b1;
    load = 1'b0;
    #1 $display("|94|%b|%b|%b|", in, load, out);

    in = 1'b1;
    load = 1'b0;
    #1 $display("|94+|%b|%b|%b|", in, load, out);

    in = 1'b1;
    load = 1'b0;
    #1 $display("|95|%b|%b|%b|", in, load, out);

    in = 1'b1;
    load = 1'b0;
    #1 $display("|95+|%b|%b|%b|", in, load, out);

    in = 1'b1;
    load = 1'b0;
    #1 $display("|96|%b|%b|%b|", in, load, out);

    in = 1'b1;
    load = 1'b0;
    #1 $display("|96+|%b|%b|%b|", in, load, out);

    in = 1'b1;
    load = 1'b0;
    #1 $display("|97|%b|%b|%b|", in, load, out);

    in = 1'b1;
    load = 1'b0;
    #1 $display("|97+|%b|%b|%b|", in, load, out);

    in = 1'b1;
    load = 1'b0;
    #1 $display("|98|%b|%b|%b|", in, load, out);

    in = 1'b1;
    load = 1'b0;
    #1 $display("|98+|%b|%b|%b|", in, load, out);

    in = 1'b1;
    load = 1'b0;
    #1 $display("|99|%b|%b|%b|", in, load, out);

    in = 1'b1;
    load = 1'b0;
    #1 $display("|99+|%b|%b|%b|", in, load, out);

    in = 1'b1;
    load = 1'b0;
    #1 $display("|100|%b|%b|%b|", in, load, out);

    in = 1'b1;
    load = 1'b0;
    #1 $display("|100+|%b|%b|%b|", in, load, out);

    in = 1'b1;
    load = 1'b0;
    #1 $display("|101|%b|%b|%b|", in, load, out);

    in = 1'b1;
    load = 1'b0;
    #1 $display("|101+|%b|%b|%b|", in, load, out);

    in = 1'b1;
    load = 1'b0;
    #1 $display("|102|%b|%b|%b|", in, load, out);

    in = 1'b1;
    load = 1'b0;
    #1 $display("|102+|%b|%b|%b|", in, load, out);

    in = 1'b1;
    load = 1'b0;
    #1 $display("|103|%b|%b|%b|", in, load, out);

    in = 1'b1;
    load = 1'b0;
    #1 $display("|103+|%b|%b|%b|", in, load, out);

    in = 1'b1;
    load = 1'b0;
    #1 $display("|104|%b|%b|%b|", in, load, out);

    in = 1'b1;
    load = 1'b0;
    #1 $display("|104+|%b|%b|%b|", in, load, out);

    in = 1'b1;
    load = 1'b0;
    #1 $display("|105|%b|%b|%b|", in, load, out);

    in = 1'b1;
    load = 1'b0;
    #1 $display("|105+|%b|%b|%b|", in, load, out);

    in = 1'b1;
    load = 1'b0;
    #1 $display("|106|%b|%b|%b|", in, load, out);

    in = 1'b1;
    load = 1'b0;
    #1 $display("|106+|%b|%b|%b|", in, load, out);

    in = 1'b1;
    load = 1'b0;
    #1 $display("|107|%b|%b|%b|", in, load, out);

    $finish;
  end
endmodule
