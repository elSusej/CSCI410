module ram64_test;
  reg signed [15:0] in;
  reg load;
  reg [5:0] address;
  wire signed [15:0] out;

  student_ram64 dut (.in(in), .load(load), .address(address), .out(out));

  initial begin
    $display("|time|in|load|address|out|");

    in = 0;
    load = 1'b0;
    address = 0;
    #1 $display("|0+|%d|%b|%d|%d|", in, load, address, out);

    in = 0;
    load = 1'b0;
    address = 0;
    #1 $display("|1|%d|%b|%d|%d|", in, load, address, out);

    in = 0;
    load = 1'b1;
    address = 0;
    #1 $display("|1+|%d|%b|%d|%d|", in, load, address, out);

    in = 0;
    load = 1'b1;
    address = 0;
    #1 $display("|2|%d|%b|%d|%d|", in, load, address, out);

    in = 1313;
    load = 1'b0;
    address = 0;
    #1 $display("|2+|%d|%b|%d|%d|", in, load, address, out);

    in = 1313;
    load = 1'b0;
    address = 0;
    #1 $display("|3|%d|%b|%d|%d|", in, load, address, out);

    in = 1313;
    load = 1'b1;
    address = 13;
    #1 $display("|3+|%d|%b|%d|%d|", in, load, address, out);

    in = 1313;
    load = 1'b1;
    address = 13;
    #1 $display("|4|%d|%b|%d|%d|", in, load, address, out);

    in = 1313;
    load = 1'b0;
    address = 0;
    #1 $display("|4+|%d|%b|%d|%d|", in, load, address, out);

    in = 1313;
    load = 1'b0;
    address = 0;
    #1 $display("|5|%d|%b|%d|%d|", in, load, address, out);

    in = 4747;
    load = 1'b0;
    address = 47;
    #1 $display("|5+|%d|%b|%d|%d|", in, load, address, out);

    in = 4747;
    load = 1'b0;
    address = 47;
    #1 $display("|6|%d|%b|%d|%d|", in, load, address, out);

    in = 4747;
    load = 1'b1;
    address = 47;
    #1 $display("|6+|%d|%b|%d|%d|", in, load, address, out);

    in = 4747;
    load = 1'b1;
    address = 47;
    #1 $display("|7|%d|%b|%d|%d|", in, load, address, out);

    in = 4747;
    load = 1'b0;
    address = 47;
    #1 $display("|7+|%d|%b|%d|%d|", in, load, address, out);

    in = 4747;
    load = 1'b0;
    address = 47;
    #1 $display("|8|%d|%b|%d|%d|", in, load, address, out);

    in = 4747;
    load = 1'b0;
    address = 13;
    #0 $display("|8|%d|%b|%d|%d|", in, load, address, out);

    in = 6363;
    load = 1'b0;
    address = 13;
    #1 $display("|8+|%d|%b|%d|%d|", in, load, address, out);

    in = 6363;
    load = 1'b0;
    address = 13;
    #1 $display("|9|%d|%b|%d|%d|", in, load, address, out);

    in = 6363;
    load = 1'b1;
    address = 63;
    #1 $display("|9+|%d|%b|%d|%d|", in, load, address, out);

    in = 6363;
    load = 1'b1;
    address = 63;
    #1 $display("|10|%d|%b|%d|%d|", in, load, address, out);

    in = 6363;
    load = 1'b0;
    address = 63;
    #1 $display("|10+|%d|%b|%d|%d|", in, load, address, out);

    in = 6363;
    load = 1'b0;
    address = 63;
    #1 $display("|11|%d|%b|%d|%d|", in, load, address, out);

    in = 6363;
    load = 1'b0;
    address = 47;
    #0 $display("|11|%d|%b|%d|%d|", in, load, address, out);

    in = 6363;
    load = 1'b0;
    address = 63;
    #0 $display("|11|%d|%b|%d|%d|", in, load, address, out);

    in = 6363;
    load = 1'b0;
    address = 40;
    #1 $display("|11+|%d|%b|%d|%d|", in, load, address, out);

    in = 6363;
    load = 1'b0;
    address = 40;
    #1 $display("|12|%d|%b|%d|%d|", in, load, address, out);

    in = 6363;
    load = 1'b0;
    address = 41;
    #0 $display("|12|%d|%b|%d|%d|", in, load, address, out);

    in = 6363;
    load = 1'b0;
    address = 42;
    #0 $display("|12|%d|%b|%d|%d|", in, load, address, out);

    in = 6363;
    load = 1'b0;
    address = 43;
    #0 $display("|12|%d|%b|%d|%d|", in, load, address, out);

    in = 6363;
    load = 1'b0;
    address = 44;
    #0 $display("|12|%d|%b|%d|%d|", in, load, address, out);

    in = 6363;
    load = 1'b0;
    address = 45;
    #0 $display("|12|%d|%b|%d|%d|", in, load, address, out);

    in = 6363;
    load = 1'b0;
    address = 46;
    #0 $display("|12|%d|%b|%d|%d|", in, load, address, out);

    in = 6363;
    load = 1'b0;
    address = 47;
    #0 $display("|12|%d|%b|%d|%d|", in, load, address, out);

    in = 21845;
    load = 1'b1;
    address = 40;
    #1 $display("|12+|%d|%b|%d|%d|", in, load, address, out);

    in = 21845;
    load = 1'b1;
    address = 40;
    #1 $display("|13|%d|%b|%d|%d|", in, load, address, out);

    in = 21845;
    load = 1'b1;
    address = 41;
    #1 $display("|13+|%d|%b|%d|%d|", in, load, address, out);

    in = 21845;
    load = 1'b1;
    address = 41;
    #1 $display("|14|%d|%b|%d|%d|", in, load, address, out);

    in = 21845;
    load = 1'b1;
    address = 42;
    #1 $display("|14+|%d|%b|%d|%d|", in, load, address, out);

    in = 21845;
    load = 1'b1;
    address = 42;
    #1 $display("|15|%d|%b|%d|%d|", in, load, address, out);

    in = 21845;
    load = 1'b1;
    address = 43;
    #1 $display("|15+|%d|%b|%d|%d|", in, load, address, out);

    in = 21845;
    load = 1'b1;
    address = 43;
    #1 $display("|16|%d|%b|%d|%d|", in, load, address, out);

    in = 21845;
    load = 1'b1;
    address = 44;
    #1 $display("|16+|%d|%b|%d|%d|", in, load, address, out);

    in = 21845;
    load = 1'b1;
    address = 44;
    #1 $display("|17|%d|%b|%d|%d|", in, load, address, out);

    in = 21845;
    load = 1'b1;
    address = 45;
    #1 $display("|17+|%d|%b|%d|%d|", in, load, address, out);

    in = 21845;
    load = 1'b1;
    address = 45;
    #1 $display("|18|%d|%b|%d|%d|", in, load, address, out);

    in = 21845;
    load = 1'b1;
    address = 46;
    #1 $display("|18+|%d|%b|%d|%d|", in, load, address, out);

    in = 21845;
    load = 1'b1;
    address = 46;
    #1 $display("|19|%d|%b|%d|%d|", in, load, address, out);

    in = 21845;
    load = 1'b1;
    address = 47;
    #1 $display("|19+|%d|%b|%d|%d|", in, load, address, out);

    in = 21845;
    load = 1'b1;
    address = 47;
    #1 $display("|20|%d|%b|%d|%d|", in, load, address, out);

    in = 21845;
    load = 1'b0;
    address = 40;
    #1 $display("|20+|%d|%b|%d|%d|", in, load, address, out);

    in = 21845;
    load = 1'b0;
    address = 40;
    #1 $display("|21|%d|%b|%d|%d|", in, load, address, out);

    in = 21845;
    load = 1'b0;
    address = 41;
    #0 $display("|21|%d|%b|%d|%d|", in, load, address, out);

    in = 21845;
    load = 1'b0;
    address = 42;
    #0 $display("|21|%d|%b|%d|%d|", in, load, address, out);

    in = 21845;
    load = 1'b0;
    address = 43;
    #0 $display("|21|%d|%b|%d|%d|", in, load, address, out);

    in = 21845;
    load = 1'b0;
    address = 44;
    #0 $display("|21|%d|%b|%d|%d|", in, load, address, out);

    in = 21845;
    load = 1'b0;
    address = 45;
    #0 $display("|21|%d|%b|%d|%d|", in, load, address, out);

    in = 21845;
    load = 1'b0;
    address = 46;
    #0 $display("|21|%d|%b|%d|%d|", in, load, address, out);

    in = 21845;
    load = 1'b0;
    address = 47;
    #0 $display("|21|%d|%b|%d|%d|", in, load, address, out);

    in = -21846;
    load = 1'b1;
    address = 40;
    #1 $display("|21+|%d|%b|%d|%d|", in, load, address, out);

    in = -21846;
    load = 1'b1;
    address = 40;
    #1 $display("|22|%d|%b|%d|%d|", in, load, address, out);

    in = -21846;
    load = 1'b0;
    address = 40;
    #1 $display("|22+|%d|%b|%d|%d|", in, load, address, out);

    in = -21846;
    load = 1'b0;
    address = 40;
    #1 $display("|23|%d|%b|%d|%d|", in, load, address, out);

    in = -21846;
    load = 1'b0;
    address = 41;
    #0 $display("|23|%d|%b|%d|%d|", in, load, address, out);

    in = -21846;
    load = 1'b0;
    address = 42;
    #0 $display("|23|%d|%b|%d|%d|", in, load, address, out);

    in = -21846;
    load = 1'b0;
    address = 43;
    #0 $display("|23|%d|%b|%d|%d|", in, load, address, out);

    in = -21846;
    load = 1'b0;
    address = 44;
    #0 $display("|23|%d|%b|%d|%d|", in, load, address, out);

    in = -21846;
    load = 1'b0;
    address = 45;
    #0 $display("|23|%d|%b|%d|%d|", in, load, address, out);

    in = -21846;
    load = 1'b0;
    address = 46;
    #0 $display("|23|%d|%b|%d|%d|", in, load, address, out);

    in = -21846;
    load = 1'b0;
    address = 47;
    #0 $display("|23|%d|%b|%d|%d|", in, load, address, out);

    in = 21845;
    load = 1'b1;
    address = 40;
    #1 $display("|23+|%d|%b|%d|%d|", in, load, address, out);

    in = 21845;
    load = 1'b1;
    address = 40;
    #1 $display("|24|%d|%b|%d|%d|", in, load, address, out);

    in = -21846;
    load = 1'b1;
    address = 41;
    #1 $display("|24+|%d|%b|%d|%d|", in, load, address, out);

    in = -21846;
    load = 1'b1;
    address = 41;
    #1 $display("|25|%d|%b|%d|%d|", in, load, address, out);

    in = -21846;
    load = 1'b0;
    address = 40;
    #1 $display("|25+|%d|%b|%d|%d|", in, load, address, out);

    in = -21846;
    load = 1'b0;
    address = 40;
    #1 $display("|26|%d|%b|%d|%d|", in, load, address, out);

    in = -21846;
    load = 1'b0;
    address = 41;
    #0 $display("|26|%d|%b|%d|%d|", in, load, address, out);

    in = -21846;
    load = 1'b0;
    address = 42;
    #0 $display("|26|%d|%b|%d|%d|", in, load, address, out);

    in = -21846;
    load = 1'b0;
    address = 43;
    #0 $display("|26|%d|%b|%d|%d|", in, load, address, out);

    in = -21846;
    load = 1'b0;
    address = 44;
    #0 $display("|26|%d|%b|%d|%d|", in, load, address, out);

    in = -21846;
    load = 1'b0;
    address = 45;
    #0 $display("|26|%d|%b|%d|%d|", in, load, address, out);

    in = -21846;
    load = 1'b0;
    address = 46;
    #0 $display("|26|%d|%b|%d|%d|", in, load, address, out);

    in = -21846;
    load = 1'b0;
    address = 47;
    #0 $display("|26|%d|%b|%d|%d|", in, load, address, out);

    in = 21845;
    load = 1'b1;
    address = 41;
    #1 $display("|26+|%d|%b|%d|%d|", in, load, address, out);

    in = 21845;
    load = 1'b1;
    address = 41;
    #1 $display("|27|%d|%b|%d|%d|", in, load, address, out);

    in = -21846;
    load = 1'b1;
    address = 42;
    #1 $display("|27+|%d|%b|%d|%d|", in, load, address, out);

    in = -21846;
    load = 1'b1;
    address = 42;
    #1 $display("|28|%d|%b|%d|%d|", in, load, address, out);

    in = -21846;
    load = 1'b0;
    address = 40;
    #1 $display("|28+|%d|%b|%d|%d|", in, load, address, out);

    in = -21846;
    load = 1'b0;
    address = 40;
    #1 $display("|29|%d|%b|%d|%d|", in, load, address, out);

    in = -21846;
    load = 1'b0;
    address = 41;
    #0 $display("|29|%d|%b|%d|%d|", in, load, address, out);

    in = -21846;
    load = 1'b0;
    address = 42;
    #0 $display("|29|%d|%b|%d|%d|", in, load, address, out);

    in = -21846;
    load = 1'b0;
    address = 43;
    #0 $display("|29|%d|%b|%d|%d|", in, load, address, out);

    in = -21846;
    load = 1'b0;
    address = 44;
    #0 $display("|29|%d|%b|%d|%d|", in, load, address, out);

    in = -21846;
    load = 1'b0;
    address = 45;
    #0 $display("|29|%d|%b|%d|%d|", in, load, address, out);

    in = -21846;
    load = 1'b0;
    address = 46;
    #0 $display("|29|%d|%b|%d|%d|", in, load, address, out);

    in = -21846;
    load = 1'b0;
    address = 47;
    #0 $display("|29|%d|%b|%d|%d|", in, load, address, out);

    in = 21845;
    load = 1'b1;
    address = 42;
    #1 $display("|29+|%d|%b|%d|%d|", in, load, address, out);

    in = 21845;
    load = 1'b1;
    address = 42;
    #1 $display("|30|%d|%b|%d|%d|", in, load, address, out);

    in = -21846;
    load = 1'b1;
    address = 43;
    #1 $display("|30+|%d|%b|%d|%d|", in, load, address, out);

    in = -21846;
    load = 1'b1;
    address = 43;
    #1 $display("|31|%d|%b|%d|%d|", in, load, address, out);

    in = -21846;
    load = 1'b0;
    address = 40;
    #1 $display("|31+|%d|%b|%d|%d|", in, load, address, out);

    in = -21846;
    load = 1'b0;
    address = 40;
    #1 $display("|32|%d|%b|%d|%d|", in, load, address, out);

    in = -21846;
    load = 1'b0;
    address = 41;
    #0 $display("|32|%d|%b|%d|%d|", in, load, address, out);

    in = -21846;
    load = 1'b0;
    address = 42;
    #0 $display("|32|%d|%b|%d|%d|", in, load, address, out);

    in = -21846;
    load = 1'b0;
    address = 43;
    #0 $display("|32|%d|%b|%d|%d|", in, load, address, out);

    in = -21846;
    load = 1'b0;
    address = 44;
    #0 $display("|32|%d|%b|%d|%d|", in, load, address, out);

    in = -21846;
    load = 1'b0;
    address = 45;
    #0 $display("|32|%d|%b|%d|%d|", in, load, address, out);

    in = -21846;
    load = 1'b0;
    address = 46;
    #0 $display("|32|%d|%b|%d|%d|", in, load, address, out);

    in = -21846;
    load = 1'b0;
    address = 47;
    #0 $display("|32|%d|%b|%d|%d|", in, load, address, out);

    in = 21845;
    load = 1'b1;
    address = 43;
    #1 $display("|32+|%d|%b|%d|%d|", in, load, address, out);

    in = 21845;
    load = 1'b1;
    address = 43;
    #1 $display("|33|%d|%b|%d|%d|", in, load, address, out);

    in = -21846;
    load = 1'b1;
    address = 44;
    #1 $display("|33+|%d|%b|%d|%d|", in, load, address, out);

    in = -21846;
    load = 1'b1;
    address = 44;
    #1 $display("|34|%d|%b|%d|%d|", in, load, address, out);

    in = -21846;
    load = 1'b0;
    address = 40;
    #1 $display("|34+|%d|%b|%d|%d|", in, load, address, out);

    in = -21846;
    load = 1'b0;
    address = 40;
    #1 $display("|35|%d|%b|%d|%d|", in, load, address, out);

    in = -21846;
    load = 1'b0;
    address = 41;
    #0 $display("|35|%d|%b|%d|%d|", in, load, address, out);

    in = -21846;
    load = 1'b0;
    address = 42;
    #0 $display("|35|%d|%b|%d|%d|", in, load, address, out);

    in = -21846;
    load = 1'b0;
    address = 43;
    #0 $display("|35|%d|%b|%d|%d|", in, load, address, out);

    in = -21846;
    load = 1'b0;
    address = 44;
    #0 $display("|35|%d|%b|%d|%d|", in, load, address, out);

    in = -21846;
    load = 1'b0;
    address = 45;
    #0 $display("|35|%d|%b|%d|%d|", in, load, address, out);

    in = -21846;
    load = 1'b0;
    address = 46;
    #0 $display("|35|%d|%b|%d|%d|", in, load, address, out);

    in = -21846;
    load = 1'b0;
    address = 47;
    #0 $display("|35|%d|%b|%d|%d|", in, load, address, out);

    in = 21845;
    load = 1'b1;
    address = 44;
    #1 $display("|35+|%d|%b|%d|%d|", in, load, address, out);

    in = 21845;
    load = 1'b1;
    address = 44;
    #1 $display("|36|%d|%b|%d|%d|", in, load, address, out);

    in = -21846;
    load = 1'b1;
    address = 45;
    #1 $display("|36+|%d|%b|%d|%d|", in, load, address, out);

    in = -21846;
    load = 1'b1;
    address = 45;
    #1 $display("|37|%d|%b|%d|%d|", in, load, address, out);

    in = -21846;
    load = 1'b0;
    address = 40;
    #1 $display("|37+|%d|%b|%d|%d|", in, load, address, out);

    in = -21846;
    load = 1'b0;
    address = 40;
    #1 $display("|38|%d|%b|%d|%d|", in, load, address, out);

    in = -21846;
    load = 1'b0;
    address = 41;
    #0 $display("|38|%d|%b|%d|%d|", in, load, address, out);

    in = -21846;
    load = 1'b0;
    address = 42;
    #0 $display("|38|%d|%b|%d|%d|", in, load, address, out);

    in = -21846;
    load = 1'b0;
    address = 43;
    #0 $display("|38|%d|%b|%d|%d|", in, load, address, out);

    in = -21846;
    load = 1'b0;
    address = 44;
    #0 $display("|38|%d|%b|%d|%d|", in, load, address, out);

    in = -21846;
    load = 1'b0;
    address = 45;
    #0 $display("|38|%d|%b|%d|%d|", in, load, address, out);

    in = -21846;
    load = 1'b0;
    address = 46;
    #0 $display("|38|%d|%b|%d|%d|", in, load, address, out);

    in = -21846;
    load = 1'b0;
    address = 47;
    #0 $display("|38|%d|%b|%d|%d|", in, load, address, out);

    in = 21845;
    load = 1'b1;
    address = 45;
    #1 $display("|38+|%d|%b|%d|%d|", in, load, address, out);

    in = 21845;
    load = 1'b1;
    address = 45;
    #1 $display("|39|%d|%b|%d|%d|", in, load, address, out);

    in = -21846;
    load = 1'b1;
    address = 46;
    #1 $display("|39+|%d|%b|%d|%d|", in, load, address, out);

    in = -21846;
    load = 1'b1;
    address = 46;
    #1 $display("|40|%d|%b|%d|%d|", in, load, address, out);

    in = -21846;
    load = 1'b0;
    address = 40;
    #1 $display("|40+|%d|%b|%d|%d|", in, load, address, out);

    in = -21846;
    load = 1'b0;
    address = 40;
    #1 $display("|41|%d|%b|%d|%d|", in, load, address, out);

    in = -21846;
    load = 1'b0;
    address = 41;
    #0 $display("|41|%d|%b|%d|%d|", in, load, address, out);

    in = -21846;
    load = 1'b0;
    address = 42;
    #0 $display("|41|%d|%b|%d|%d|", in, load, address, out);

    in = -21846;
    load = 1'b0;
    address = 43;
    #0 $display("|41|%d|%b|%d|%d|", in, load, address, out);

    in = -21846;
    load = 1'b0;
    address = 44;
    #0 $display("|41|%d|%b|%d|%d|", in, load, address, out);

    in = -21846;
    load = 1'b0;
    address = 45;
    #0 $display("|41|%d|%b|%d|%d|", in, load, address, out);

    in = -21846;
    load = 1'b0;
    address = 46;
    #0 $display("|41|%d|%b|%d|%d|", in, load, address, out);

    in = -21846;
    load = 1'b0;
    address = 47;
    #0 $display("|41|%d|%b|%d|%d|", in, load, address, out);

    in = 21845;
    load = 1'b1;
    address = 46;
    #1 $display("|41+|%d|%b|%d|%d|", in, load, address, out);

    in = 21845;
    load = 1'b1;
    address = 46;
    #1 $display("|42|%d|%b|%d|%d|", in, load, address, out);

    in = -21846;
    load = 1'b1;
    address = 47;
    #1 $display("|42+|%d|%b|%d|%d|", in, load, address, out);

    in = -21846;
    load = 1'b1;
    address = 47;
    #1 $display("|43|%d|%b|%d|%d|", in, load, address, out);

    in = -21846;
    load = 1'b0;
    address = 40;
    #1 $display("|43+|%d|%b|%d|%d|", in, load, address, out);

    in = -21846;
    load = 1'b0;
    address = 40;
    #1 $display("|44|%d|%b|%d|%d|", in, load, address, out);

    in = -21846;
    load = 1'b0;
    address = 41;
    #0 $display("|44|%d|%b|%d|%d|", in, load, address, out);

    in = -21846;
    load = 1'b0;
    address = 42;
    #0 $display("|44|%d|%b|%d|%d|", in, load, address, out);

    in = -21846;
    load = 1'b0;
    address = 43;
    #0 $display("|44|%d|%b|%d|%d|", in, load, address, out);

    in = -21846;
    load = 1'b0;
    address = 44;
    #0 $display("|44|%d|%b|%d|%d|", in, load, address, out);

    in = -21846;
    load = 1'b0;
    address = 45;
    #0 $display("|44|%d|%b|%d|%d|", in, load, address, out);

    in = -21846;
    load = 1'b0;
    address = 46;
    #0 $display("|44|%d|%b|%d|%d|", in, load, address, out);

    in = -21846;
    load = 1'b0;
    address = 47;
    #0 $display("|44|%d|%b|%d|%d|", in, load, address, out);

    in = 21845;
    load = 1'b1;
    address = 47;
    #1 $display("|44+|%d|%b|%d|%d|", in, load, address, out);

    in = 21845;
    load = 1'b1;
    address = 47;
    #1 $display("|45|%d|%b|%d|%d|", in, load, address, out);

    in = 21845;
    load = 1'b0;
    address = 40;
    #1 $display("|45+|%d|%b|%d|%d|", in, load, address, out);

    in = 21845;
    load = 1'b0;
    address = 40;
    #1 $display("|46|%d|%b|%d|%d|", in, load, address, out);

    in = 21845;
    load = 1'b0;
    address = 41;
    #0 $display("|46|%d|%b|%d|%d|", in, load, address, out);

    in = 21845;
    load = 1'b0;
    address = 42;
    #0 $display("|46|%d|%b|%d|%d|", in, load, address, out);

    in = 21845;
    load = 1'b0;
    address = 43;
    #0 $display("|46|%d|%b|%d|%d|", in, load, address, out);

    in = 21845;
    load = 1'b0;
    address = 44;
    #0 $display("|46|%d|%b|%d|%d|", in, load, address, out);

    in = 21845;
    load = 1'b0;
    address = 45;
    #0 $display("|46|%d|%b|%d|%d|", in, load, address, out);

    in = 21845;
    load = 1'b0;
    address = 46;
    #0 $display("|46|%d|%b|%d|%d|", in, load, address, out);

    in = 21845;
    load = 1'b0;
    address = 47;
    #0 $display("|46|%d|%b|%d|%d|", in, load, address, out);

    in = 21845;
    load = 1'b0;
    address = 5;
    #1 $display("|46+|%d|%b|%d|%d|", in, load, address, out);

    in = 21845;
    load = 1'b0;
    address = 5;
    #1 $display("|47|%d|%b|%d|%d|", in, load, address, out);

    in = 21845;
    load = 1'b0;
    address = 13;
    #0 $display("|47|%d|%b|%d|%d|", in, load, address, out);

    in = 21845;
    load = 1'b0;
    address = 21;
    #0 $display("|47|%d|%b|%d|%d|", in, load, address, out);

    in = 21845;
    load = 1'b0;
    address = 29;
    #0 $display("|47|%d|%b|%d|%d|", in, load, address, out);

    in = 21845;
    load = 1'b0;
    address = 37;
    #0 $display("|47|%d|%b|%d|%d|", in, load, address, out);

    in = 21845;
    load = 1'b0;
    address = 45;
    #0 $display("|47|%d|%b|%d|%d|", in, load, address, out);

    in = 21845;
    load = 1'b0;
    address = 53;
    #0 $display("|47|%d|%b|%d|%d|", in, load, address, out);

    in = 21845;
    load = 1'b0;
    address = 61;
    #0 $display("|47|%d|%b|%d|%d|", in, load, address, out);

    in = 21845;
    load = 1'b1;
    address = 5;
    #1 $display("|47+|%d|%b|%d|%d|", in, load, address, out);

    in = 21845;
    load = 1'b1;
    address = 5;
    #1 $display("|48|%d|%b|%d|%d|", in, load, address, out);

    in = 21845;
    load = 1'b1;
    address = 13;
    #1 $display("|48+|%d|%b|%d|%d|", in, load, address, out);

    in = 21845;
    load = 1'b1;
    address = 13;
    #1 $display("|49|%d|%b|%d|%d|", in, load, address, out);

    in = 21845;
    load = 1'b1;
    address = 21;
    #1 $display("|49+|%d|%b|%d|%d|", in, load, address, out);

    in = 21845;
    load = 1'b1;
    address = 21;
    #1 $display("|50|%d|%b|%d|%d|", in, load, address, out);

    in = 21845;
    load = 1'b1;
    address = 29;
    #1 $display("|50+|%d|%b|%d|%d|", in, load, address, out);

    in = 21845;
    load = 1'b1;
    address = 29;
    #1 $display("|51|%d|%b|%d|%d|", in, load, address, out);

    in = 21845;
    load = 1'b1;
    address = 37;
    #1 $display("|51+|%d|%b|%d|%d|", in, load, address, out);

    in = 21845;
    load = 1'b1;
    address = 37;
    #1 $display("|52|%d|%b|%d|%d|", in, load, address, out);

    in = 21845;
    load = 1'b1;
    address = 45;
    #1 $display("|52+|%d|%b|%d|%d|", in, load, address, out);

    in = 21845;
    load = 1'b1;
    address = 45;
    #1 $display("|53|%d|%b|%d|%d|", in, load, address, out);

    in = 21845;
    load = 1'b1;
    address = 53;
    #1 $display("|53+|%d|%b|%d|%d|", in, load, address, out);

    in = 21845;
    load = 1'b1;
    address = 53;
    #1 $display("|54|%d|%b|%d|%d|", in, load, address, out);

    in = 21845;
    load = 1'b1;
    address = 61;
    #1 $display("|54+|%d|%b|%d|%d|", in, load, address, out);

    in = 21845;
    load = 1'b1;
    address = 61;
    #1 $display("|55|%d|%b|%d|%d|", in, load, address, out);

    in = 21845;
    load = 1'b0;
    address = 5;
    #1 $display("|55+|%d|%b|%d|%d|", in, load, address, out);

    in = 21845;
    load = 1'b0;
    address = 5;
    #1 $display("|56|%d|%b|%d|%d|", in, load, address, out);

    in = 21845;
    load = 1'b0;
    address = 13;
    #0 $display("|56|%d|%b|%d|%d|", in, load, address, out);

    in = 21845;
    load = 1'b0;
    address = 21;
    #0 $display("|56|%d|%b|%d|%d|", in, load, address, out);

    in = 21845;
    load = 1'b0;
    address = 29;
    #0 $display("|56|%d|%b|%d|%d|", in, load, address, out);

    in = 21845;
    load = 1'b0;
    address = 37;
    #0 $display("|56|%d|%b|%d|%d|", in, load, address, out);

    in = 21845;
    load = 1'b0;
    address = 45;
    #0 $display("|56|%d|%b|%d|%d|", in, load, address, out);

    in = 21845;
    load = 1'b0;
    address = 53;
    #0 $display("|56|%d|%b|%d|%d|", in, load, address, out);

    in = 21845;
    load = 1'b0;
    address = 61;
    #0 $display("|56|%d|%b|%d|%d|", in, load, address, out);

    in = -21846;
    load = 1'b1;
    address = 5;
    #1 $display("|56+|%d|%b|%d|%d|", in, load, address, out);

    in = -21846;
    load = 1'b1;
    address = 5;
    #1 $display("|57|%d|%b|%d|%d|", in, load, address, out);

    in = -21846;
    load = 1'b0;
    address = 5;
    #1 $display("|57+|%d|%b|%d|%d|", in, load, address, out);

    in = -21846;
    load = 1'b0;
    address = 5;
    #1 $display("|58|%d|%b|%d|%d|", in, load, address, out);

    in = -21846;
    load = 1'b0;
    address = 13;
    #0 $display("|58|%d|%b|%d|%d|", in, load, address, out);

    in = -21846;
    load = 1'b0;
    address = 21;
    #0 $display("|58|%d|%b|%d|%d|", in, load, address, out);

    in = -21846;
    load = 1'b0;
    address = 29;
    #0 $display("|58|%d|%b|%d|%d|", in, load, address, out);

    in = -21846;
    load = 1'b0;
    address = 37;
    #0 $display("|58|%d|%b|%d|%d|", in, load, address, out);

    in = -21846;
    load = 1'b0;
    address = 45;
    #0 $display("|58|%d|%b|%d|%d|", in, load, address, out);

    in = -21846;
    load = 1'b0;
    address = 53;
    #0 $display("|58|%d|%b|%d|%d|", in, load, address, out);

    in = -21846;
    load = 1'b0;
    address = 61;
    #0 $display("|58|%d|%b|%d|%d|", in, load, address, out);

    in = 21845;
    load = 1'b1;
    address = 5;
    #1 $display("|58+|%d|%b|%d|%d|", in, load, address, out);

    in = 21845;
    load = 1'b1;
    address = 5;
    #1 $display("|59|%d|%b|%d|%d|", in, load, address, out);

    in = -21846;
    load = 1'b1;
    address = 13;
    #1 $display("|59+|%d|%b|%d|%d|", in, load, address, out);

    in = -21846;
    load = 1'b1;
    address = 13;
    #1 $display("|60|%d|%b|%d|%d|", in, load, address, out);

    in = -21846;
    load = 1'b0;
    address = 5;
    #1 $display("|60+|%d|%b|%d|%d|", in, load, address, out);

    in = -21846;
    load = 1'b0;
    address = 5;
    #1 $display("|61|%d|%b|%d|%d|", in, load, address, out);

    in = -21846;
    load = 1'b0;
    address = 13;
    #0 $display("|61|%d|%b|%d|%d|", in, load, address, out);

    in = -21846;
    load = 1'b0;
    address = 21;
    #0 $display("|61|%d|%b|%d|%d|", in, load, address, out);

    in = -21846;
    load = 1'b0;
    address = 29;
    #0 $display("|61|%d|%b|%d|%d|", in, load, address, out);

    in = -21846;
    load = 1'b0;
    address = 37;
    #0 $display("|61|%d|%b|%d|%d|", in, load, address, out);

    in = -21846;
    load = 1'b0;
    address = 45;
    #0 $display("|61|%d|%b|%d|%d|", in, load, address, out);

    in = -21846;
    load = 1'b0;
    address = 53;
    #0 $display("|61|%d|%b|%d|%d|", in, load, address, out);

    in = -21846;
    load = 1'b0;
    address = 61;
    #0 $display("|61|%d|%b|%d|%d|", in, load, address, out);

    in = 21845;
    load = 1'b1;
    address = 13;
    #1 $display("|61+|%d|%b|%d|%d|", in, load, address, out);

    in = 21845;
    load = 1'b1;
    address = 13;
    #1 $display("|62|%d|%b|%d|%d|", in, load, address, out);

    in = -21846;
    load = 1'b1;
    address = 21;
    #1 $display("|62+|%d|%b|%d|%d|", in, load, address, out);

    in = -21846;
    load = 1'b1;
    address = 21;
    #1 $display("|63|%d|%b|%d|%d|", in, load, address, out);

    in = -21846;
    load = 1'b0;
    address = 5;
    #1 $display("|63+|%d|%b|%d|%d|", in, load, address, out);

    in = -21846;
    load = 1'b0;
    address = 5;
    #1 $display("|64|%d|%b|%d|%d|", in, load, address, out);

    in = -21846;
    load = 1'b0;
    address = 13;
    #0 $display("|64|%d|%b|%d|%d|", in, load, address, out);

    in = -21846;
    load = 1'b0;
    address = 21;
    #0 $display("|64|%d|%b|%d|%d|", in, load, address, out);

    in = -21846;
    load = 1'b0;
    address = 29;
    #0 $display("|64|%d|%b|%d|%d|", in, load, address, out);

    in = -21846;
    load = 1'b0;
    address = 37;
    #0 $display("|64|%d|%b|%d|%d|", in, load, address, out);

    in = -21846;
    load = 1'b0;
    address = 45;
    #0 $display("|64|%d|%b|%d|%d|", in, load, address, out);

    in = -21846;
    load = 1'b0;
    address = 53;
    #0 $display("|64|%d|%b|%d|%d|", in, load, address, out);

    in = -21846;
    load = 1'b0;
    address = 61;
    #0 $display("|64|%d|%b|%d|%d|", in, load, address, out);

    in = 21845;
    load = 1'b1;
    address = 21;
    #1 $display("|64+|%d|%b|%d|%d|", in, load, address, out);

    in = 21845;
    load = 1'b1;
    address = 21;
    #1 $display("|65|%d|%b|%d|%d|", in, load, address, out);

    in = -21846;
    load = 1'b1;
    address = 29;
    #1 $display("|65+|%d|%b|%d|%d|", in, load, address, out);

    in = -21846;
    load = 1'b1;
    address = 29;
    #1 $display("|66|%d|%b|%d|%d|", in, load, address, out);

    in = -21846;
    load = 1'b0;
    address = 5;
    #1 $display("|66+|%d|%b|%d|%d|", in, load, address, out);

    in = -21846;
    load = 1'b0;
    address = 5;
    #1 $display("|67|%d|%b|%d|%d|", in, load, address, out);

    in = -21846;
    load = 1'b0;
    address = 13;
    #0 $display("|67|%d|%b|%d|%d|", in, load, address, out);

    in = -21846;
    load = 1'b0;
    address = 21;
    #0 $display("|67|%d|%b|%d|%d|", in, load, address, out);

    in = -21846;
    load = 1'b0;
    address = 29;
    #0 $display("|67|%d|%b|%d|%d|", in, load, address, out);

    in = -21846;
    load = 1'b0;
    address = 37;
    #0 $display("|67|%d|%b|%d|%d|", in, load, address, out);

    in = -21846;
    load = 1'b0;
    address = 45;
    #0 $display("|67|%d|%b|%d|%d|", in, load, address, out);

    in = -21846;
    load = 1'b0;
    address = 53;
    #0 $display("|67|%d|%b|%d|%d|", in, load, address, out);

    in = -21846;
    load = 1'b0;
    address = 61;
    #0 $display("|67|%d|%b|%d|%d|", in, load, address, out);

    in = 21845;
    load = 1'b1;
    address = 29;
    #1 $display("|67+|%d|%b|%d|%d|", in, load, address, out);

    in = 21845;
    load = 1'b1;
    address = 29;
    #1 $display("|68|%d|%b|%d|%d|", in, load, address, out);

    in = -21846;
    load = 1'b1;
    address = 37;
    #1 $display("|68+|%d|%b|%d|%d|", in, load, address, out);

    in = -21846;
    load = 1'b1;
    address = 37;
    #1 $display("|69|%d|%b|%d|%d|", in, load, address, out);

    in = -21846;
    load = 1'b0;
    address = 5;
    #1 $display("|69+|%d|%b|%d|%d|", in, load, address, out);

    in = -21846;
    load = 1'b0;
    address = 5;
    #1 $display("|70|%d|%b|%d|%d|", in, load, address, out);

    in = -21846;
    load = 1'b0;
    address = 13;
    #0 $display("|70|%d|%b|%d|%d|", in, load, address, out);

    in = -21846;
    load = 1'b0;
    address = 21;
    #0 $display("|70|%d|%b|%d|%d|", in, load, address, out);

    in = -21846;
    load = 1'b0;
    address = 29;
    #0 $display("|70|%d|%b|%d|%d|", in, load, address, out);

    in = -21846;
    load = 1'b0;
    address = 37;
    #0 $display("|70|%d|%b|%d|%d|", in, load, address, out);

    in = -21846;
    load = 1'b0;
    address = 45;
    #0 $display("|70|%d|%b|%d|%d|", in, load, address, out);

    in = -21846;
    load = 1'b0;
    address = 53;
    #0 $display("|70|%d|%b|%d|%d|", in, load, address, out);

    in = -21846;
    load = 1'b0;
    address = 61;
    #0 $display("|70|%d|%b|%d|%d|", in, load, address, out);

    in = 21845;
    load = 1'b1;
    address = 37;
    #1 $display("|70+|%d|%b|%d|%d|", in, load, address, out);

    in = 21845;
    load = 1'b1;
    address = 37;
    #1 $display("|71|%d|%b|%d|%d|", in, load, address, out);

    in = -21846;
    load = 1'b1;
    address = 45;
    #1 $display("|71+|%d|%b|%d|%d|", in, load, address, out);

    in = -21846;
    load = 1'b1;
    address = 45;
    #1 $display("|72|%d|%b|%d|%d|", in, load, address, out);

    in = -21846;
    load = 1'b0;
    address = 5;
    #1 $display("|72+|%d|%b|%d|%d|", in, load, address, out);

    in = -21846;
    load = 1'b0;
    address = 5;
    #1 $display("|73|%d|%b|%d|%d|", in, load, address, out);

    in = -21846;
    load = 1'b0;
    address = 13;
    #0 $display("|73|%d|%b|%d|%d|", in, load, address, out);

    in = -21846;
    load = 1'b0;
    address = 21;
    #0 $display("|73|%d|%b|%d|%d|", in, load, address, out);

    in = -21846;
    load = 1'b0;
    address = 29;
    #0 $display("|73|%d|%b|%d|%d|", in, load, address, out);

    in = -21846;
    load = 1'b0;
    address = 37;
    #0 $display("|73|%d|%b|%d|%d|", in, load, address, out);

    in = -21846;
    load = 1'b0;
    address = 45;
    #0 $display("|73|%d|%b|%d|%d|", in, load, address, out);

    in = -21846;
    load = 1'b0;
    address = 53;
    #0 $display("|73|%d|%b|%d|%d|", in, load, address, out);

    in = -21846;
    load = 1'b0;
    address = 61;
    #0 $display("|73|%d|%b|%d|%d|", in, load, address, out);

    in = 21845;
    load = 1'b1;
    address = 45;
    #1 $display("|73+|%d|%b|%d|%d|", in, load, address, out);

    in = 21845;
    load = 1'b1;
    address = 45;
    #1 $display("|74|%d|%b|%d|%d|", in, load, address, out);

    in = -21846;
    load = 1'b1;
    address = 53;
    #1 $display("|74+|%d|%b|%d|%d|", in, load, address, out);

    in = -21846;
    load = 1'b1;
    address = 53;
    #1 $display("|75|%d|%b|%d|%d|", in, load, address, out);

    in = -21846;
    load = 1'b0;
    address = 5;
    #1 $display("|75+|%d|%b|%d|%d|", in, load, address, out);

    in = -21846;
    load = 1'b0;
    address = 5;
    #1 $display("|76|%d|%b|%d|%d|", in, load, address, out);

    in = -21846;
    load = 1'b0;
    address = 13;
    #0 $display("|76|%d|%b|%d|%d|", in, load, address, out);

    in = -21846;
    load = 1'b0;
    address = 21;
    #0 $display("|76|%d|%b|%d|%d|", in, load, address, out);

    in = -21846;
    load = 1'b0;
    address = 29;
    #0 $display("|76|%d|%b|%d|%d|", in, load, address, out);

    in = -21846;
    load = 1'b0;
    address = 37;
    #0 $display("|76|%d|%b|%d|%d|", in, load, address, out);

    in = -21846;
    load = 1'b0;
    address = 45;
    #0 $display("|76|%d|%b|%d|%d|", in, load, address, out);

    in = -21846;
    load = 1'b0;
    address = 53;
    #0 $display("|76|%d|%b|%d|%d|", in, load, address, out);

    in = -21846;
    load = 1'b0;
    address = 61;
    #0 $display("|76|%d|%b|%d|%d|", in, load, address, out);

    in = 21845;
    load = 1'b1;
    address = 53;
    #1 $display("|76+|%d|%b|%d|%d|", in, load, address, out);

    in = 21845;
    load = 1'b1;
    address = 53;
    #1 $display("|77|%d|%b|%d|%d|", in, load, address, out);

    in = -21846;
    load = 1'b1;
    address = 61;
    #1 $display("|77+|%d|%b|%d|%d|", in, load, address, out);

    in = -21846;
    load = 1'b1;
    address = 61;
    #1 $display("|78|%d|%b|%d|%d|", in, load, address, out);

    in = -21846;
    load = 1'b0;
    address = 5;
    #1 $display("|78+|%d|%b|%d|%d|", in, load, address, out);

    in = -21846;
    load = 1'b0;
    address = 5;
    #1 $display("|79|%d|%b|%d|%d|", in, load, address, out);

    in = -21846;
    load = 1'b0;
    address = 13;
    #0 $display("|79|%d|%b|%d|%d|", in, load, address, out);

    in = -21846;
    load = 1'b0;
    address = 21;
    #0 $display("|79|%d|%b|%d|%d|", in, load, address, out);

    in = -21846;
    load = 1'b0;
    address = 29;
    #0 $display("|79|%d|%b|%d|%d|", in, load, address, out);

    in = -21846;
    load = 1'b0;
    address = 37;
    #0 $display("|79|%d|%b|%d|%d|", in, load, address, out);

    in = -21846;
    load = 1'b0;
    address = 45;
    #0 $display("|79|%d|%b|%d|%d|", in, load, address, out);

    in = -21846;
    load = 1'b0;
    address = 53;
    #0 $display("|79|%d|%b|%d|%d|", in, load, address, out);

    in = -21846;
    load = 1'b0;
    address = 61;
    #0 $display("|79|%d|%b|%d|%d|", in, load, address, out);

    in = 21845;
    load = 1'b1;
    address = 61;
    #1 $display("|79+|%d|%b|%d|%d|", in, load, address, out);

    in = 21845;
    load = 1'b1;
    address = 61;
    #1 $display("|80|%d|%b|%d|%d|", in, load, address, out);

    in = 21845;
    load = 1'b0;
    address = 5;
    #1 $display("|80+|%d|%b|%d|%d|", in, load, address, out);

    in = 21845;
    load = 1'b0;
    address = 5;
    #1 $display("|81|%d|%b|%d|%d|", in, load, address, out);

    in = 21845;
    load = 1'b0;
    address = 13;
    #0 $display("|81|%d|%b|%d|%d|", in, load, address, out);

    in = 21845;
    load = 1'b0;
    address = 21;
    #0 $display("|81|%d|%b|%d|%d|", in, load, address, out);

    in = 21845;
    load = 1'b0;
    address = 29;
    #0 $display("|81|%d|%b|%d|%d|", in, load, address, out);

    in = 21845;
    load = 1'b0;
    address = 37;
    #0 $display("|81|%d|%b|%d|%d|", in, load, address, out);

    in = 21845;
    load = 1'b0;
    address = 45;
    #0 $display("|81|%d|%b|%d|%d|", in, load, address, out);

    in = 21845;
    load = 1'b0;
    address = 53;
    #0 $display("|81|%d|%b|%d|%d|", in, load, address, out);

    in = 21845;
    load = 1'b0;
    address = 61;
    #0 $display("|81|%d|%b|%d|%d|", in, load, address, out);

    $finish;
  end
endmodule
